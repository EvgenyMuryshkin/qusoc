----------------------------------------------------------------------------------------------------------------------------------
-- libraries
----------------------------------------------------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all;

----------------------------------------------------------------------------------------------------------------------------------
-- entity declaration
----------------------------------------------------------------------------------------------------------------------------------
entity fir_iq_sym_decimator_ram is
    generic(
          g_outreg                  : integer := 1
        ; g_ram_size                : integer := 32
    );
    port(
          CLK                       : in std_logic
        ; CE                        : in std_logic
        ; WR                        : in std_logic
        ; WR_ADDR                   : in std_logic_vector(4 downto 0)
        ; DIN                       : in std_logic_vector(15 downto 0)
        ; RD                        : in std_logic
        ; RD_ADDR                   : in std_logic_vector(4 downto 0)
        ; DOUT                      : out std_logic_vector(15 downto 0)
    );
end entity;

----------------------------------------------------------------------------------------------------------------------------------
-- architecture declaration
----------------------------------------------------------------------------------------------------------------------------------
architecture behavioral of fir_iq_sym_decimator_ram is
	type slv16_array is array (0 to g_ram_size - 1) of std_logic_vector (15 downto 0);
----------------------------------------------------------------------------------------------------------------------------------
-- signals declaration
----------------------------------------------------------------------------------------------------------------------------------
    signal
        ib_din
            : std_logic_vector(15 downto 0) := (others => '0');
--    signal
    signal
        ram
            : slv16_array := (others => (others => '0'));

    signal
        ram_out_r1,
        ram_out_r2
            : std_logic_vector(15 downto 0) := (others => '0');

begin
----------------------------------------------------------------------------------------------------------------------------------
-- input
----------------------------------------------------------------------------------------------------------------------------------
    ib_din                          <= DIN;

----------------------------------------------------------------------------------------------------------------------------------
-- process, write/read ram
----------------------------------------------------------------------------------------------------------------------------------
    p_ram : process(CLK)
    begin
        if (rising_edge(CLK)) then
				if (CE = '1' and WR = '1') then                    
					ram(conv_integer(WR_ADDR)) <= ib_din;
				end if; -- CE

				if (CE = '1' and RD = '1') then
                    if (g_outreg = 1) then
                        ram_out_r2 <= ram(conv_integer(RD_ADDR));
                    elsif (g_outreg = 2) then
                        ram_out_r1 <= ram(conv_integer(RD_ADDR));
                        ram_out_r2 <= ram_out_r1;
                    end if;
				end if; -- CE
			              
        end if; -- CLK
    end process;

----------------------------------------------------------------------------------------------------------------------------------
-- output
----------------------------------------------------------------------------------------------------------------------------------
    DOUT                            <= ram_out_r2;

----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
end;