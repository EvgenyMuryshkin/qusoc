`timescale 1ns/1ps
`default_nettype none

`define Assert(expected, actual, message) \
if (expected !== actual) begin \
$display("Assert failed"); \
$display(message); \
$display("Expected: 0x%H, Actual: 0x%H", expected, actual); \
/*$finish;*/ \
end

module VGASyncModule_testbench;
	reg clk;
	reg reset;

	reg Enabled;

	wire OutVisible;
	wire OutFP;
	wire OutSP;
	wire OutBP;
	wire OutMax;
	wire [9:0] OutCounter;

	initial begin
		clk = 1'b0;
		forever clk = #500 ~clk;
	end

	initial begin
		reset = 1'b1;
		@(negedge clk);
		reset = 1'b0;

	end

	initial begin

		Enabled = 1'b0;
		@(negedge clk); // reset

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 1");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 1");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 1");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 1");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 1");
		`Assert(10'b0000000001, OutCounter, "OutCounter: value does not match at clock 1");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 2");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 2");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 2");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 2");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 2");
		`Assert(10'b0000000010, OutCounter, "OutCounter: value does not match at clock 2");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 3");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 3");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 3");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 3");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 3");
		`Assert(10'b0000000011, OutCounter, "OutCounter: value does not match at clock 3");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 4");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 4");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 4");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 4");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 4");
		`Assert(10'b0000000100, OutCounter, "OutCounter: value does not match at clock 4");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 5");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 5");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 5");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 5");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 5");
		`Assert(10'b0000000101, OutCounter, "OutCounter: value does not match at clock 5");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 6");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 6");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 6");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 6");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 6");
		`Assert(10'b0000000110, OutCounter, "OutCounter: value does not match at clock 6");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 7");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 7");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 7");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 7");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 7");
		`Assert(10'b0000000111, OutCounter, "OutCounter: value does not match at clock 7");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 8");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 8");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 8");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 8");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 8");
		`Assert(10'b0000001000, OutCounter, "OutCounter: value does not match at clock 8");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 9");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 9");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 9");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 9");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 9");
		`Assert(10'b0000001001, OutCounter, "OutCounter: value does not match at clock 9");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 10");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 10");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 10");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 10");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 10");
		`Assert(10'b0000001010, OutCounter, "OutCounter: value does not match at clock 10");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 11");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 11");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 11");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 11");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 11");
		`Assert(10'b0000001011, OutCounter, "OutCounter: value does not match at clock 11");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 12");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 12");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 12");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 12");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 12");
		`Assert(10'b0000001100, OutCounter, "OutCounter: value does not match at clock 12");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 13");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 13");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 13");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 13");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 13");
		`Assert(10'b0000001101, OutCounter, "OutCounter: value does not match at clock 13");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 14");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 14");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 14");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 14");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 14");
		`Assert(10'b0000001110, OutCounter, "OutCounter: value does not match at clock 14");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 15");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 15");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 15");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 15");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 15");
		`Assert(10'b0000001111, OutCounter, "OutCounter: value does not match at clock 15");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 16");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 16");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 16");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 16");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 16");
		`Assert(10'b0000010000, OutCounter, "OutCounter: value does not match at clock 16");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 17");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 17");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 17");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 17");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 17");
		`Assert(10'b0000010001, OutCounter, "OutCounter: value does not match at clock 17");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 18");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 18");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 18");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 18");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 18");
		`Assert(10'b0000010010, OutCounter, "OutCounter: value does not match at clock 18");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 19");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 19");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 19");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 19");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 19");
		`Assert(10'b0000010011, OutCounter, "OutCounter: value does not match at clock 19");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 20");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 20");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 20");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 20");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 20");
		`Assert(10'b0000010100, OutCounter, "OutCounter: value does not match at clock 20");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 21");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 21");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 21");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 21");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 21");
		`Assert(10'b0000010101, OutCounter, "OutCounter: value does not match at clock 21");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 22");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 22");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 22");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 22");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 22");
		`Assert(10'b0000010110, OutCounter, "OutCounter: value does not match at clock 22");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 23");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 23");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 23");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 23");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 23");
		`Assert(10'b0000010111, OutCounter, "OutCounter: value does not match at clock 23");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 24");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 24");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 24");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 24");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 24");
		`Assert(10'b0000011000, OutCounter, "OutCounter: value does not match at clock 24");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 25");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 25");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 25");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 25");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 25");
		`Assert(10'b0000011001, OutCounter, "OutCounter: value does not match at clock 25");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 26");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 26");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 26");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 26");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 26");
		`Assert(10'b0000011010, OutCounter, "OutCounter: value does not match at clock 26");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 27");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 27");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 27");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 27");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 27");
		`Assert(10'b0000011011, OutCounter, "OutCounter: value does not match at clock 27");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 28");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 28");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 28");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 28");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 28");
		`Assert(10'b0000011100, OutCounter, "OutCounter: value does not match at clock 28");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 29");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 29");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 29");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 29");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 29");
		`Assert(10'b0000011101, OutCounter, "OutCounter: value does not match at clock 29");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 30");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 30");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 30");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 30");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 30");
		`Assert(10'b0000011110, OutCounter, "OutCounter: value does not match at clock 30");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 31");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 31");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 31");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 31");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 31");
		`Assert(10'b0000011111, OutCounter, "OutCounter: value does not match at clock 31");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 32");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 32");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 32");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 32");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 32");
		`Assert(10'b0000100000, OutCounter, "OutCounter: value does not match at clock 32");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 33");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 33");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 33");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 33");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 33");
		`Assert(10'b0000100001, OutCounter, "OutCounter: value does not match at clock 33");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 34");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 34");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 34");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 34");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 34");
		`Assert(10'b0000100010, OutCounter, "OutCounter: value does not match at clock 34");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 35");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 35");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 35");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 35");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 35");
		`Assert(10'b0000100011, OutCounter, "OutCounter: value does not match at clock 35");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 36");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 36");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 36");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 36");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 36");
		`Assert(10'b0000100100, OutCounter, "OutCounter: value does not match at clock 36");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 37");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 37");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 37");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 37");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 37");
		`Assert(10'b0000100101, OutCounter, "OutCounter: value does not match at clock 37");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 38");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 38");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 38");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 38");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 38");
		`Assert(10'b0000100110, OutCounter, "OutCounter: value does not match at clock 38");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 39");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 39");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 39");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 39");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 39");
		`Assert(10'b0000100111, OutCounter, "OutCounter: value does not match at clock 39");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 40");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 40");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 40");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 40");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 40");
		`Assert(10'b0000101000, OutCounter, "OutCounter: value does not match at clock 40");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 41");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 41");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 41");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 41");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 41");
		`Assert(10'b0000101001, OutCounter, "OutCounter: value does not match at clock 41");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 42");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 42");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 42");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 42");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 42");
		`Assert(10'b0000101010, OutCounter, "OutCounter: value does not match at clock 42");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 43");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 43");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 43");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 43");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 43");
		`Assert(10'b0000101011, OutCounter, "OutCounter: value does not match at clock 43");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 44");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 44");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 44");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 44");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 44");
		`Assert(10'b0000101100, OutCounter, "OutCounter: value does not match at clock 44");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 45");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 45");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 45");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 45");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 45");
		`Assert(10'b0000101101, OutCounter, "OutCounter: value does not match at clock 45");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 46");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 46");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 46");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 46");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 46");
		`Assert(10'b0000101110, OutCounter, "OutCounter: value does not match at clock 46");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 47");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 47");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 47");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 47");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 47");
		`Assert(10'b0000101111, OutCounter, "OutCounter: value does not match at clock 47");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 48");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 48");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 48");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 48");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 48");
		`Assert(10'b0000110000, OutCounter, "OutCounter: value does not match at clock 48");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 49");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 49");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 49");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 49");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 49");
		`Assert(10'b0000110001, OutCounter, "OutCounter: value does not match at clock 49");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 50");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 50");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 50");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 50");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 50");
		`Assert(10'b0000110010, OutCounter, "OutCounter: value does not match at clock 50");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 51");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 51");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 51");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 51");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 51");
		`Assert(10'b0000110011, OutCounter, "OutCounter: value does not match at clock 51");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 52");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 52");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 52");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 52");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 52");
		`Assert(10'b0000110100, OutCounter, "OutCounter: value does not match at clock 52");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 53");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 53");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 53");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 53");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 53");
		`Assert(10'b0000110101, OutCounter, "OutCounter: value does not match at clock 53");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 54");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 54");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 54");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 54");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 54");
		`Assert(10'b0000110110, OutCounter, "OutCounter: value does not match at clock 54");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 55");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 55");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 55");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 55");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 55");
		`Assert(10'b0000110111, OutCounter, "OutCounter: value does not match at clock 55");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 56");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 56");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 56");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 56");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 56");
		`Assert(10'b0000111000, OutCounter, "OutCounter: value does not match at clock 56");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 57");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 57");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 57");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 57");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 57");
		`Assert(10'b0000111001, OutCounter, "OutCounter: value does not match at clock 57");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 58");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 58");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 58");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 58");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 58");
		`Assert(10'b0000111010, OutCounter, "OutCounter: value does not match at clock 58");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 59");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 59");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 59");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 59");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 59");
		`Assert(10'b0000111011, OutCounter, "OutCounter: value does not match at clock 59");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 60");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 60");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 60");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 60");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 60");
		`Assert(10'b0000111100, OutCounter, "OutCounter: value does not match at clock 60");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 61");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 61");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 61");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 61");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 61");
		`Assert(10'b0000111101, OutCounter, "OutCounter: value does not match at clock 61");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 62");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 62");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 62");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 62");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 62");
		`Assert(10'b0000111110, OutCounter, "OutCounter: value does not match at clock 62");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 63");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 63");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 63");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 63");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 63");
		`Assert(10'b0000111111, OutCounter, "OutCounter: value does not match at clock 63");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 64");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 64");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 64");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 64");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 64");
		`Assert(10'b0001000000, OutCounter, "OutCounter: value does not match at clock 64");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 65");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 65");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 65");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 65");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 65");
		`Assert(10'b0001000001, OutCounter, "OutCounter: value does not match at clock 65");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 66");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 66");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 66");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 66");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 66");
		`Assert(10'b0001000010, OutCounter, "OutCounter: value does not match at clock 66");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 67");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 67");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 67");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 67");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 67");
		`Assert(10'b0001000011, OutCounter, "OutCounter: value does not match at clock 67");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 68");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 68");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 68");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 68");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 68");
		`Assert(10'b0001000100, OutCounter, "OutCounter: value does not match at clock 68");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 69");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 69");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 69");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 69");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 69");
		`Assert(10'b0001000101, OutCounter, "OutCounter: value does not match at clock 69");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 70");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 70");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 70");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 70");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 70");
		`Assert(10'b0001000110, OutCounter, "OutCounter: value does not match at clock 70");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 71");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 71");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 71");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 71");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 71");
		`Assert(10'b0001000111, OutCounter, "OutCounter: value does not match at clock 71");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 72");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 72");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 72");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 72");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 72");
		`Assert(10'b0001001000, OutCounter, "OutCounter: value does not match at clock 72");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 73");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 73");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 73");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 73");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 73");
		`Assert(10'b0001001001, OutCounter, "OutCounter: value does not match at clock 73");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 74");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 74");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 74");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 74");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 74");
		`Assert(10'b0001001010, OutCounter, "OutCounter: value does not match at clock 74");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 75");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 75");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 75");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 75");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 75");
		`Assert(10'b0001001011, OutCounter, "OutCounter: value does not match at clock 75");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 76");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 76");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 76");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 76");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 76");
		`Assert(10'b0001001100, OutCounter, "OutCounter: value does not match at clock 76");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 77");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 77");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 77");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 77");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 77");
		`Assert(10'b0001001101, OutCounter, "OutCounter: value does not match at clock 77");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 78");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 78");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 78");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 78");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 78");
		`Assert(10'b0001001110, OutCounter, "OutCounter: value does not match at clock 78");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 79");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 79");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 79");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 79");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 79");
		`Assert(10'b0001001111, OutCounter, "OutCounter: value does not match at clock 79");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 80");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 80");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 80");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 80");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 80");
		`Assert(10'b0001010000, OutCounter, "OutCounter: value does not match at clock 80");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 81");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 81");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 81");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 81");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 81");
		`Assert(10'b0001010001, OutCounter, "OutCounter: value does not match at clock 81");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 82");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 82");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 82");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 82");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 82");
		`Assert(10'b0001010010, OutCounter, "OutCounter: value does not match at clock 82");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 83");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 83");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 83");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 83");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 83");
		`Assert(10'b0001010011, OutCounter, "OutCounter: value does not match at clock 83");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 84");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 84");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 84");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 84");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 84");
		`Assert(10'b0001010100, OutCounter, "OutCounter: value does not match at clock 84");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 85");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 85");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 85");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 85");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 85");
		`Assert(10'b0001010101, OutCounter, "OutCounter: value does not match at clock 85");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 86");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 86");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 86");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 86");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 86");
		`Assert(10'b0001010110, OutCounter, "OutCounter: value does not match at clock 86");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 87");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 87");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 87");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 87");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 87");
		`Assert(10'b0001010111, OutCounter, "OutCounter: value does not match at clock 87");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 88");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 88");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 88");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 88");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 88");
		`Assert(10'b0001011000, OutCounter, "OutCounter: value does not match at clock 88");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 89");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 89");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 89");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 89");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 89");
		`Assert(10'b0001011001, OutCounter, "OutCounter: value does not match at clock 89");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 90");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 90");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 90");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 90");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 90");
		`Assert(10'b0001011010, OutCounter, "OutCounter: value does not match at clock 90");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 91");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 91");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 91");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 91");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 91");
		`Assert(10'b0001011011, OutCounter, "OutCounter: value does not match at clock 91");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 92");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 92");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 92");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 92");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 92");
		`Assert(10'b0001011100, OutCounter, "OutCounter: value does not match at clock 92");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 93");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 93");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 93");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 93");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 93");
		`Assert(10'b0001011101, OutCounter, "OutCounter: value does not match at clock 93");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 94");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 94");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 94");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 94");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 94");
		`Assert(10'b0001011110, OutCounter, "OutCounter: value does not match at clock 94");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 95");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 95");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 95");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 95");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 95");
		`Assert(10'b0001011111, OutCounter, "OutCounter: value does not match at clock 95");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 96");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 96");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 96");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 96");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 96");
		`Assert(10'b0001100000, OutCounter, "OutCounter: value does not match at clock 96");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 97");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 97");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 97");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 97");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 97");
		`Assert(10'b0001100001, OutCounter, "OutCounter: value does not match at clock 97");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 98");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 98");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 98");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 98");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 98");
		`Assert(10'b0001100010, OutCounter, "OutCounter: value does not match at clock 98");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 99");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 99");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 99");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 99");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 99");
		`Assert(10'b0001100011, OutCounter, "OutCounter: value does not match at clock 99");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 100");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 100");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 100");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 100");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 100");
		`Assert(10'b0001100100, OutCounter, "OutCounter: value does not match at clock 100");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 101");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 101");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 101");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 101");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 101");
		`Assert(10'b0001100101, OutCounter, "OutCounter: value does not match at clock 101");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 102");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 102");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 102");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 102");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 102");
		`Assert(10'b0001100110, OutCounter, "OutCounter: value does not match at clock 102");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 103");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 103");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 103");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 103");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 103");
		`Assert(10'b0001100111, OutCounter, "OutCounter: value does not match at clock 103");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 104");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 104");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 104");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 104");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 104");
		`Assert(10'b0001101000, OutCounter, "OutCounter: value does not match at clock 104");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 105");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 105");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 105");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 105");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 105");
		`Assert(10'b0001101001, OutCounter, "OutCounter: value does not match at clock 105");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 106");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 106");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 106");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 106");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 106");
		`Assert(10'b0001101010, OutCounter, "OutCounter: value does not match at clock 106");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 107");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 107");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 107");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 107");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 107");
		`Assert(10'b0001101011, OutCounter, "OutCounter: value does not match at clock 107");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 108");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 108");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 108");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 108");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 108");
		`Assert(10'b0001101100, OutCounter, "OutCounter: value does not match at clock 108");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 109");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 109");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 109");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 109");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 109");
		`Assert(10'b0001101101, OutCounter, "OutCounter: value does not match at clock 109");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 110");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 110");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 110");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 110");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 110");
		`Assert(10'b0001101110, OutCounter, "OutCounter: value does not match at clock 110");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 111");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 111");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 111");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 111");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 111");
		`Assert(10'b0001101111, OutCounter, "OutCounter: value does not match at clock 111");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 112");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 112");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 112");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 112");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 112");
		`Assert(10'b0001110000, OutCounter, "OutCounter: value does not match at clock 112");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 113");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 113");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 113");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 113");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 113");
		`Assert(10'b0001110001, OutCounter, "OutCounter: value does not match at clock 113");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 114");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 114");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 114");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 114");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 114");
		`Assert(10'b0001110010, OutCounter, "OutCounter: value does not match at clock 114");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 115");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 115");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 115");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 115");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 115");
		`Assert(10'b0001110011, OutCounter, "OutCounter: value does not match at clock 115");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 116");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 116");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 116");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 116");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 116");
		`Assert(10'b0001110100, OutCounter, "OutCounter: value does not match at clock 116");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 117");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 117");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 117");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 117");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 117");
		`Assert(10'b0001110101, OutCounter, "OutCounter: value does not match at clock 117");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 118");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 118");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 118");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 118");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 118");
		`Assert(10'b0001110110, OutCounter, "OutCounter: value does not match at clock 118");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 119");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 119");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 119");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 119");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 119");
		`Assert(10'b0001110111, OutCounter, "OutCounter: value does not match at clock 119");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 120");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 120");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 120");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 120");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 120");
		`Assert(10'b0001111000, OutCounter, "OutCounter: value does not match at clock 120");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 121");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 121");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 121");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 121");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 121");
		`Assert(10'b0001111001, OutCounter, "OutCounter: value does not match at clock 121");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 122");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 122");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 122");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 122");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 122");
		`Assert(10'b0001111010, OutCounter, "OutCounter: value does not match at clock 122");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 123");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 123");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 123");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 123");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 123");
		`Assert(10'b0001111011, OutCounter, "OutCounter: value does not match at clock 123");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 124");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 124");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 124");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 124");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 124");
		`Assert(10'b0001111100, OutCounter, "OutCounter: value does not match at clock 124");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 125");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 125");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 125");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 125");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 125");
		`Assert(10'b0001111101, OutCounter, "OutCounter: value does not match at clock 125");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 126");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 126");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 126");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 126");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 126");
		`Assert(10'b0001111110, OutCounter, "OutCounter: value does not match at clock 126");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 127");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 127");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 127");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 127");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 127");
		`Assert(10'b0001111111, OutCounter, "OutCounter: value does not match at clock 127");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 128");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 128");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 128");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 128");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 128");
		`Assert(10'b0010000000, OutCounter, "OutCounter: value does not match at clock 128");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 129");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 129");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 129");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 129");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 129");
		`Assert(10'b0010000001, OutCounter, "OutCounter: value does not match at clock 129");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 130");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 130");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 130");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 130");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 130");
		`Assert(10'b0010000010, OutCounter, "OutCounter: value does not match at clock 130");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 131");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 131");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 131");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 131");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 131");
		`Assert(10'b0010000011, OutCounter, "OutCounter: value does not match at clock 131");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 132");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 132");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 132");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 132");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 132");
		`Assert(10'b0010000100, OutCounter, "OutCounter: value does not match at clock 132");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 133");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 133");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 133");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 133");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 133");
		`Assert(10'b0010000101, OutCounter, "OutCounter: value does not match at clock 133");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 134");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 134");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 134");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 134");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 134");
		`Assert(10'b0010000110, OutCounter, "OutCounter: value does not match at clock 134");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 135");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 135");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 135");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 135");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 135");
		`Assert(10'b0010000111, OutCounter, "OutCounter: value does not match at clock 135");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 136");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 136");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 136");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 136");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 136");
		`Assert(10'b0010001000, OutCounter, "OutCounter: value does not match at clock 136");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 137");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 137");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 137");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 137");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 137");
		`Assert(10'b0010001001, OutCounter, "OutCounter: value does not match at clock 137");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 138");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 138");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 138");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 138");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 138");
		`Assert(10'b0010001010, OutCounter, "OutCounter: value does not match at clock 138");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 139");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 139");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 139");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 139");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 139");
		`Assert(10'b0010001011, OutCounter, "OutCounter: value does not match at clock 139");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 140");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 140");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 140");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 140");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 140");
		`Assert(10'b0010001100, OutCounter, "OutCounter: value does not match at clock 140");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 141");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 141");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 141");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 141");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 141");
		`Assert(10'b0010001101, OutCounter, "OutCounter: value does not match at clock 141");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 142");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 142");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 142");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 142");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 142");
		`Assert(10'b0010001110, OutCounter, "OutCounter: value does not match at clock 142");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 143");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 143");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 143");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 143");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 143");
		`Assert(10'b0010001111, OutCounter, "OutCounter: value does not match at clock 143");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 144");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 144");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 144");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 144");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 144");
		`Assert(10'b0010010000, OutCounter, "OutCounter: value does not match at clock 144");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 145");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 145");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 145");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 145");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 145");
		`Assert(10'b0010010001, OutCounter, "OutCounter: value does not match at clock 145");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 146");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 146");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 146");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 146");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 146");
		`Assert(10'b0010010010, OutCounter, "OutCounter: value does not match at clock 146");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 147");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 147");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 147");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 147");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 147");
		`Assert(10'b0010010011, OutCounter, "OutCounter: value does not match at clock 147");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 148");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 148");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 148");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 148");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 148");
		`Assert(10'b0010010100, OutCounter, "OutCounter: value does not match at clock 148");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 149");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 149");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 149");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 149");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 149");
		`Assert(10'b0010010101, OutCounter, "OutCounter: value does not match at clock 149");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 150");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 150");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 150");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 150");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 150");
		`Assert(10'b0010010110, OutCounter, "OutCounter: value does not match at clock 150");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 151");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 151");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 151");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 151");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 151");
		`Assert(10'b0010010111, OutCounter, "OutCounter: value does not match at clock 151");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 152");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 152");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 152");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 152");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 152");
		`Assert(10'b0010011000, OutCounter, "OutCounter: value does not match at clock 152");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 153");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 153");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 153");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 153");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 153");
		`Assert(10'b0010011001, OutCounter, "OutCounter: value does not match at clock 153");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 154");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 154");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 154");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 154");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 154");
		`Assert(10'b0010011010, OutCounter, "OutCounter: value does not match at clock 154");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 155");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 155");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 155");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 155");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 155");
		`Assert(10'b0010011011, OutCounter, "OutCounter: value does not match at clock 155");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 156");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 156");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 156");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 156");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 156");
		`Assert(10'b0010011100, OutCounter, "OutCounter: value does not match at clock 156");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 157");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 157");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 157");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 157");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 157");
		`Assert(10'b0010011101, OutCounter, "OutCounter: value does not match at clock 157");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 158");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 158");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 158");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 158");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 158");
		`Assert(10'b0010011110, OutCounter, "OutCounter: value does not match at clock 158");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 159");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 159");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 159");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 159");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 159");
		`Assert(10'b0010011111, OutCounter, "OutCounter: value does not match at clock 159");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 160");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 160");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 160");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 160");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 160");
		`Assert(10'b0010100000, OutCounter, "OutCounter: value does not match at clock 160");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 161");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 161");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 161");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 161");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 161");
		`Assert(10'b0010100001, OutCounter, "OutCounter: value does not match at clock 161");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 162");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 162");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 162");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 162");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 162");
		`Assert(10'b0010100010, OutCounter, "OutCounter: value does not match at clock 162");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 163");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 163");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 163");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 163");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 163");
		`Assert(10'b0010100011, OutCounter, "OutCounter: value does not match at clock 163");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 164");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 164");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 164");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 164");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 164");
		`Assert(10'b0010100100, OutCounter, "OutCounter: value does not match at clock 164");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 165");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 165");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 165");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 165");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 165");
		`Assert(10'b0010100101, OutCounter, "OutCounter: value does not match at clock 165");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 166");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 166");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 166");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 166");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 166");
		`Assert(10'b0010100110, OutCounter, "OutCounter: value does not match at clock 166");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 167");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 167");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 167");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 167");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 167");
		`Assert(10'b0010100111, OutCounter, "OutCounter: value does not match at clock 167");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 168");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 168");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 168");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 168");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 168");
		`Assert(10'b0010101000, OutCounter, "OutCounter: value does not match at clock 168");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 169");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 169");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 169");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 169");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 169");
		`Assert(10'b0010101001, OutCounter, "OutCounter: value does not match at clock 169");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 170");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 170");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 170");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 170");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 170");
		`Assert(10'b0010101010, OutCounter, "OutCounter: value does not match at clock 170");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 171");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 171");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 171");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 171");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 171");
		`Assert(10'b0010101011, OutCounter, "OutCounter: value does not match at clock 171");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 172");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 172");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 172");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 172");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 172");
		`Assert(10'b0010101100, OutCounter, "OutCounter: value does not match at clock 172");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 173");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 173");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 173");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 173");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 173");
		`Assert(10'b0010101101, OutCounter, "OutCounter: value does not match at clock 173");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 174");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 174");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 174");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 174");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 174");
		`Assert(10'b0010101110, OutCounter, "OutCounter: value does not match at clock 174");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 175");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 175");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 175");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 175");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 175");
		`Assert(10'b0010101111, OutCounter, "OutCounter: value does not match at clock 175");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 176");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 176");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 176");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 176");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 176");
		`Assert(10'b0010110000, OutCounter, "OutCounter: value does not match at clock 176");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 177");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 177");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 177");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 177");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 177");
		`Assert(10'b0010110001, OutCounter, "OutCounter: value does not match at clock 177");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 178");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 178");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 178");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 178");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 178");
		`Assert(10'b0010110010, OutCounter, "OutCounter: value does not match at clock 178");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 179");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 179");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 179");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 179");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 179");
		`Assert(10'b0010110011, OutCounter, "OutCounter: value does not match at clock 179");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 180");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 180");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 180");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 180");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 180");
		`Assert(10'b0010110100, OutCounter, "OutCounter: value does not match at clock 180");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 181");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 181");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 181");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 181");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 181");
		`Assert(10'b0010110101, OutCounter, "OutCounter: value does not match at clock 181");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 182");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 182");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 182");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 182");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 182");
		`Assert(10'b0010110110, OutCounter, "OutCounter: value does not match at clock 182");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 183");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 183");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 183");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 183");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 183");
		`Assert(10'b0010110111, OutCounter, "OutCounter: value does not match at clock 183");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 184");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 184");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 184");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 184");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 184");
		`Assert(10'b0010111000, OutCounter, "OutCounter: value does not match at clock 184");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 185");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 185");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 185");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 185");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 185");
		`Assert(10'b0010111001, OutCounter, "OutCounter: value does not match at clock 185");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 186");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 186");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 186");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 186");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 186");
		`Assert(10'b0010111010, OutCounter, "OutCounter: value does not match at clock 186");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 187");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 187");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 187");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 187");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 187");
		`Assert(10'b0010111011, OutCounter, "OutCounter: value does not match at clock 187");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 188");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 188");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 188");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 188");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 188");
		`Assert(10'b0010111100, OutCounter, "OutCounter: value does not match at clock 188");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 189");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 189");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 189");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 189");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 189");
		`Assert(10'b0010111101, OutCounter, "OutCounter: value does not match at clock 189");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 190");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 190");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 190");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 190");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 190");
		`Assert(10'b0010111110, OutCounter, "OutCounter: value does not match at clock 190");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 191");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 191");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 191");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 191");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 191");
		`Assert(10'b0010111111, OutCounter, "OutCounter: value does not match at clock 191");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 192");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 192");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 192");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 192");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 192");
		`Assert(10'b0011000000, OutCounter, "OutCounter: value does not match at clock 192");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 193");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 193");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 193");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 193");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 193");
		`Assert(10'b0011000001, OutCounter, "OutCounter: value does not match at clock 193");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 194");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 194");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 194");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 194");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 194");
		`Assert(10'b0011000010, OutCounter, "OutCounter: value does not match at clock 194");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 195");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 195");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 195");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 195");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 195");
		`Assert(10'b0011000011, OutCounter, "OutCounter: value does not match at clock 195");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 196");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 196");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 196");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 196");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 196");
		`Assert(10'b0011000100, OutCounter, "OutCounter: value does not match at clock 196");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 197");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 197");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 197");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 197");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 197");
		`Assert(10'b0011000101, OutCounter, "OutCounter: value does not match at clock 197");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 198");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 198");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 198");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 198");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 198");
		`Assert(10'b0011000110, OutCounter, "OutCounter: value does not match at clock 198");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 199");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 199");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 199");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 199");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 199");
		`Assert(10'b0011000111, OutCounter, "OutCounter: value does not match at clock 199");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 200");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 200");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 200");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 200");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 200");
		`Assert(10'b0011001000, OutCounter, "OutCounter: value does not match at clock 200");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 201");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 201");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 201");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 201");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 201");
		`Assert(10'b0011001001, OutCounter, "OutCounter: value does not match at clock 201");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 202");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 202");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 202");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 202");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 202");
		`Assert(10'b0011001010, OutCounter, "OutCounter: value does not match at clock 202");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 203");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 203");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 203");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 203");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 203");
		`Assert(10'b0011001011, OutCounter, "OutCounter: value does not match at clock 203");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 204");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 204");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 204");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 204");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 204");
		`Assert(10'b0011001100, OutCounter, "OutCounter: value does not match at clock 204");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 205");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 205");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 205");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 205");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 205");
		`Assert(10'b0011001101, OutCounter, "OutCounter: value does not match at clock 205");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 206");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 206");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 206");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 206");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 206");
		`Assert(10'b0011001110, OutCounter, "OutCounter: value does not match at clock 206");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 207");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 207");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 207");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 207");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 207");
		`Assert(10'b0011001111, OutCounter, "OutCounter: value does not match at clock 207");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 208");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 208");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 208");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 208");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 208");
		`Assert(10'b0011010000, OutCounter, "OutCounter: value does not match at clock 208");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 209");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 209");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 209");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 209");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 209");
		`Assert(10'b0011010001, OutCounter, "OutCounter: value does not match at clock 209");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 210");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 210");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 210");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 210");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 210");
		`Assert(10'b0011010010, OutCounter, "OutCounter: value does not match at clock 210");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 211");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 211");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 211");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 211");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 211");
		`Assert(10'b0011010011, OutCounter, "OutCounter: value does not match at clock 211");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 212");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 212");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 212");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 212");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 212");
		`Assert(10'b0011010100, OutCounter, "OutCounter: value does not match at clock 212");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 213");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 213");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 213");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 213");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 213");
		`Assert(10'b0011010101, OutCounter, "OutCounter: value does not match at clock 213");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 214");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 214");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 214");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 214");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 214");
		`Assert(10'b0011010110, OutCounter, "OutCounter: value does not match at clock 214");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 215");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 215");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 215");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 215");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 215");
		`Assert(10'b0011010111, OutCounter, "OutCounter: value does not match at clock 215");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 216");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 216");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 216");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 216");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 216");
		`Assert(10'b0011011000, OutCounter, "OutCounter: value does not match at clock 216");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 217");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 217");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 217");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 217");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 217");
		`Assert(10'b0011011001, OutCounter, "OutCounter: value does not match at clock 217");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 218");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 218");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 218");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 218");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 218");
		`Assert(10'b0011011010, OutCounter, "OutCounter: value does not match at clock 218");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 219");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 219");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 219");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 219");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 219");
		`Assert(10'b0011011011, OutCounter, "OutCounter: value does not match at clock 219");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 220");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 220");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 220");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 220");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 220");
		`Assert(10'b0011011100, OutCounter, "OutCounter: value does not match at clock 220");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 221");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 221");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 221");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 221");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 221");
		`Assert(10'b0011011101, OutCounter, "OutCounter: value does not match at clock 221");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 222");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 222");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 222");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 222");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 222");
		`Assert(10'b0011011110, OutCounter, "OutCounter: value does not match at clock 222");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 223");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 223");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 223");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 223");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 223");
		`Assert(10'b0011011111, OutCounter, "OutCounter: value does not match at clock 223");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 224");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 224");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 224");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 224");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 224");
		`Assert(10'b0011100000, OutCounter, "OutCounter: value does not match at clock 224");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 225");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 225");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 225");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 225");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 225");
		`Assert(10'b0011100001, OutCounter, "OutCounter: value does not match at clock 225");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 226");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 226");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 226");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 226");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 226");
		`Assert(10'b0011100010, OutCounter, "OutCounter: value does not match at clock 226");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 227");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 227");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 227");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 227");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 227");
		`Assert(10'b0011100011, OutCounter, "OutCounter: value does not match at clock 227");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 228");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 228");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 228");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 228");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 228");
		`Assert(10'b0011100100, OutCounter, "OutCounter: value does not match at clock 228");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 229");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 229");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 229");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 229");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 229");
		`Assert(10'b0011100101, OutCounter, "OutCounter: value does not match at clock 229");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 230");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 230");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 230");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 230");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 230");
		`Assert(10'b0011100110, OutCounter, "OutCounter: value does not match at clock 230");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 231");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 231");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 231");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 231");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 231");
		`Assert(10'b0011100111, OutCounter, "OutCounter: value does not match at clock 231");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 232");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 232");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 232");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 232");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 232");
		`Assert(10'b0011101000, OutCounter, "OutCounter: value does not match at clock 232");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 233");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 233");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 233");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 233");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 233");
		`Assert(10'b0011101001, OutCounter, "OutCounter: value does not match at clock 233");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 234");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 234");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 234");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 234");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 234");
		`Assert(10'b0011101010, OutCounter, "OutCounter: value does not match at clock 234");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 235");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 235");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 235");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 235");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 235");
		`Assert(10'b0011101011, OutCounter, "OutCounter: value does not match at clock 235");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 236");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 236");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 236");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 236");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 236");
		`Assert(10'b0011101100, OutCounter, "OutCounter: value does not match at clock 236");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 237");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 237");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 237");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 237");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 237");
		`Assert(10'b0011101101, OutCounter, "OutCounter: value does not match at clock 237");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 238");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 238");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 238");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 238");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 238");
		`Assert(10'b0011101110, OutCounter, "OutCounter: value does not match at clock 238");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 239");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 239");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 239");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 239");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 239");
		`Assert(10'b0011101111, OutCounter, "OutCounter: value does not match at clock 239");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 240");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 240");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 240");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 240");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 240");
		`Assert(10'b0011110000, OutCounter, "OutCounter: value does not match at clock 240");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 241");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 241");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 241");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 241");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 241");
		`Assert(10'b0011110001, OutCounter, "OutCounter: value does not match at clock 241");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 242");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 242");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 242");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 242");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 242");
		`Assert(10'b0011110010, OutCounter, "OutCounter: value does not match at clock 242");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 243");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 243");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 243");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 243");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 243");
		`Assert(10'b0011110011, OutCounter, "OutCounter: value does not match at clock 243");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 244");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 244");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 244");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 244");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 244");
		`Assert(10'b0011110100, OutCounter, "OutCounter: value does not match at clock 244");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 245");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 245");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 245");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 245");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 245");
		`Assert(10'b0011110101, OutCounter, "OutCounter: value does not match at clock 245");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 246");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 246");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 246");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 246");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 246");
		`Assert(10'b0011110110, OutCounter, "OutCounter: value does not match at clock 246");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 247");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 247");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 247");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 247");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 247");
		`Assert(10'b0011110111, OutCounter, "OutCounter: value does not match at clock 247");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 248");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 248");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 248");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 248");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 248");
		`Assert(10'b0011111000, OutCounter, "OutCounter: value does not match at clock 248");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 249");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 249");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 249");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 249");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 249");
		`Assert(10'b0011111001, OutCounter, "OutCounter: value does not match at clock 249");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 250");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 250");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 250");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 250");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 250");
		`Assert(10'b0011111010, OutCounter, "OutCounter: value does not match at clock 250");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 251");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 251");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 251");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 251");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 251");
		`Assert(10'b0011111011, OutCounter, "OutCounter: value does not match at clock 251");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 252");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 252");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 252");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 252");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 252");
		`Assert(10'b0011111100, OutCounter, "OutCounter: value does not match at clock 252");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 253");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 253");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 253");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 253");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 253");
		`Assert(10'b0011111101, OutCounter, "OutCounter: value does not match at clock 253");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 254");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 254");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 254");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 254");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 254");
		`Assert(10'b0011111110, OutCounter, "OutCounter: value does not match at clock 254");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 255");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 255");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 255");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 255");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 255");
		`Assert(10'b0011111111, OutCounter, "OutCounter: value does not match at clock 255");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 256");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 256");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 256");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 256");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 256");
		`Assert(10'b0100000000, OutCounter, "OutCounter: value does not match at clock 256");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 257");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 257");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 257");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 257");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 257");
		`Assert(10'b0100000001, OutCounter, "OutCounter: value does not match at clock 257");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 258");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 258");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 258");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 258");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 258");
		`Assert(10'b0100000010, OutCounter, "OutCounter: value does not match at clock 258");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 259");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 259");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 259");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 259");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 259");
		`Assert(10'b0100000011, OutCounter, "OutCounter: value does not match at clock 259");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 260");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 260");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 260");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 260");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 260");
		`Assert(10'b0100000100, OutCounter, "OutCounter: value does not match at clock 260");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 261");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 261");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 261");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 261");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 261");
		`Assert(10'b0100000101, OutCounter, "OutCounter: value does not match at clock 261");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 262");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 262");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 262");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 262");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 262");
		`Assert(10'b0100000110, OutCounter, "OutCounter: value does not match at clock 262");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 263");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 263");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 263");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 263");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 263");
		`Assert(10'b0100000111, OutCounter, "OutCounter: value does not match at clock 263");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 264");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 264");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 264");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 264");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 264");
		`Assert(10'b0100001000, OutCounter, "OutCounter: value does not match at clock 264");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 265");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 265");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 265");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 265");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 265");
		`Assert(10'b0100001001, OutCounter, "OutCounter: value does not match at clock 265");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 266");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 266");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 266");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 266");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 266");
		`Assert(10'b0100001010, OutCounter, "OutCounter: value does not match at clock 266");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 267");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 267");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 267");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 267");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 267");
		`Assert(10'b0100001011, OutCounter, "OutCounter: value does not match at clock 267");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 268");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 268");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 268");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 268");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 268");
		`Assert(10'b0100001100, OutCounter, "OutCounter: value does not match at clock 268");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 269");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 269");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 269");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 269");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 269");
		`Assert(10'b0100001101, OutCounter, "OutCounter: value does not match at clock 269");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 270");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 270");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 270");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 270");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 270");
		`Assert(10'b0100001110, OutCounter, "OutCounter: value does not match at clock 270");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 271");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 271");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 271");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 271");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 271");
		`Assert(10'b0100001111, OutCounter, "OutCounter: value does not match at clock 271");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 272");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 272");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 272");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 272");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 272");
		`Assert(10'b0100010000, OutCounter, "OutCounter: value does not match at clock 272");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 273");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 273");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 273");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 273");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 273");
		`Assert(10'b0100010001, OutCounter, "OutCounter: value does not match at clock 273");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 274");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 274");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 274");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 274");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 274");
		`Assert(10'b0100010010, OutCounter, "OutCounter: value does not match at clock 274");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 275");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 275");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 275");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 275");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 275");
		`Assert(10'b0100010011, OutCounter, "OutCounter: value does not match at clock 275");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 276");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 276");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 276");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 276");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 276");
		`Assert(10'b0100010100, OutCounter, "OutCounter: value does not match at clock 276");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 277");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 277");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 277");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 277");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 277");
		`Assert(10'b0100010101, OutCounter, "OutCounter: value does not match at clock 277");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 278");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 278");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 278");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 278");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 278");
		`Assert(10'b0100010110, OutCounter, "OutCounter: value does not match at clock 278");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 279");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 279");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 279");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 279");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 279");
		`Assert(10'b0100010111, OutCounter, "OutCounter: value does not match at clock 279");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 280");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 280");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 280");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 280");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 280");
		`Assert(10'b0100011000, OutCounter, "OutCounter: value does not match at clock 280");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 281");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 281");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 281");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 281");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 281");
		`Assert(10'b0100011001, OutCounter, "OutCounter: value does not match at clock 281");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 282");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 282");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 282");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 282");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 282");
		`Assert(10'b0100011010, OutCounter, "OutCounter: value does not match at clock 282");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 283");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 283");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 283");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 283");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 283");
		`Assert(10'b0100011011, OutCounter, "OutCounter: value does not match at clock 283");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 284");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 284");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 284");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 284");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 284");
		`Assert(10'b0100011100, OutCounter, "OutCounter: value does not match at clock 284");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 285");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 285");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 285");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 285");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 285");
		`Assert(10'b0100011101, OutCounter, "OutCounter: value does not match at clock 285");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 286");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 286");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 286");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 286");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 286");
		`Assert(10'b0100011110, OutCounter, "OutCounter: value does not match at clock 286");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 287");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 287");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 287");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 287");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 287");
		`Assert(10'b0100011111, OutCounter, "OutCounter: value does not match at clock 287");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 288");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 288");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 288");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 288");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 288");
		`Assert(10'b0100100000, OutCounter, "OutCounter: value does not match at clock 288");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 289");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 289");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 289");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 289");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 289");
		`Assert(10'b0100100001, OutCounter, "OutCounter: value does not match at clock 289");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 290");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 290");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 290");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 290");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 290");
		`Assert(10'b0100100010, OutCounter, "OutCounter: value does not match at clock 290");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 291");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 291");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 291");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 291");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 291");
		`Assert(10'b0100100011, OutCounter, "OutCounter: value does not match at clock 291");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 292");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 292");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 292");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 292");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 292");
		`Assert(10'b0100100100, OutCounter, "OutCounter: value does not match at clock 292");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 293");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 293");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 293");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 293");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 293");
		`Assert(10'b0100100101, OutCounter, "OutCounter: value does not match at clock 293");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 294");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 294");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 294");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 294");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 294");
		`Assert(10'b0100100110, OutCounter, "OutCounter: value does not match at clock 294");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 295");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 295");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 295");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 295");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 295");
		`Assert(10'b0100100111, OutCounter, "OutCounter: value does not match at clock 295");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 296");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 296");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 296");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 296");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 296");
		`Assert(10'b0100101000, OutCounter, "OutCounter: value does not match at clock 296");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 297");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 297");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 297");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 297");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 297");
		`Assert(10'b0100101001, OutCounter, "OutCounter: value does not match at clock 297");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 298");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 298");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 298");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 298");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 298");
		`Assert(10'b0100101010, OutCounter, "OutCounter: value does not match at clock 298");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 299");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 299");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 299");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 299");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 299");
		`Assert(10'b0100101011, OutCounter, "OutCounter: value does not match at clock 299");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 300");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 300");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 300");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 300");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 300");
		`Assert(10'b0100101100, OutCounter, "OutCounter: value does not match at clock 300");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 301");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 301");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 301");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 301");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 301");
		`Assert(10'b0100101101, OutCounter, "OutCounter: value does not match at clock 301");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 302");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 302");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 302");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 302");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 302");
		`Assert(10'b0100101110, OutCounter, "OutCounter: value does not match at clock 302");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 303");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 303");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 303");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 303");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 303");
		`Assert(10'b0100101111, OutCounter, "OutCounter: value does not match at clock 303");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 304");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 304");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 304");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 304");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 304");
		`Assert(10'b0100110000, OutCounter, "OutCounter: value does not match at clock 304");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 305");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 305");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 305");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 305");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 305");
		`Assert(10'b0100110001, OutCounter, "OutCounter: value does not match at clock 305");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 306");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 306");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 306");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 306");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 306");
		`Assert(10'b0100110010, OutCounter, "OutCounter: value does not match at clock 306");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 307");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 307");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 307");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 307");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 307");
		`Assert(10'b0100110011, OutCounter, "OutCounter: value does not match at clock 307");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 308");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 308");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 308");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 308");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 308");
		`Assert(10'b0100110100, OutCounter, "OutCounter: value does not match at clock 308");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 309");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 309");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 309");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 309");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 309");
		`Assert(10'b0100110101, OutCounter, "OutCounter: value does not match at clock 309");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 310");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 310");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 310");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 310");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 310");
		`Assert(10'b0100110110, OutCounter, "OutCounter: value does not match at clock 310");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 311");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 311");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 311");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 311");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 311");
		`Assert(10'b0100110111, OutCounter, "OutCounter: value does not match at clock 311");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 312");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 312");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 312");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 312");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 312");
		`Assert(10'b0100111000, OutCounter, "OutCounter: value does not match at clock 312");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 313");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 313");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 313");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 313");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 313");
		`Assert(10'b0100111001, OutCounter, "OutCounter: value does not match at clock 313");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 314");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 314");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 314");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 314");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 314");
		`Assert(10'b0100111010, OutCounter, "OutCounter: value does not match at clock 314");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 315");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 315");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 315");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 315");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 315");
		`Assert(10'b0100111011, OutCounter, "OutCounter: value does not match at clock 315");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 316");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 316");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 316");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 316");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 316");
		`Assert(10'b0100111100, OutCounter, "OutCounter: value does not match at clock 316");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 317");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 317");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 317");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 317");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 317");
		`Assert(10'b0100111101, OutCounter, "OutCounter: value does not match at clock 317");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 318");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 318");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 318");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 318");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 318");
		`Assert(10'b0100111110, OutCounter, "OutCounter: value does not match at clock 318");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 319");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 319");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 319");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 319");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 319");
		`Assert(10'b0100111111, OutCounter, "OutCounter: value does not match at clock 319");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 320");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 320");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 320");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 320");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 320");
		`Assert(10'b0101000000, OutCounter, "OutCounter: value does not match at clock 320");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 321");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 321");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 321");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 321");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 321");
		`Assert(10'b0101000001, OutCounter, "OutCounter: value does not match at clock 321");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 322");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 322");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 322");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 322");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 322");
		`Assert(10'b0101000010, OutCounter, "OutCounter: value does not match at clock 322");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 323");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 323");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 323");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 323");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 323");
		`Assert(10'b0101000011, OutCounter, "OutCounter: value does not match at clock 323");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 324");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 324");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 324");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 324");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 324");
		`Assert(10'b0101000100, OutCounter, "OutCounter: value does not match at clock 324");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 325");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 325");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 325");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 325");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 325");
		`Assert(10'b0101000101, OutCounter, "OutCounter: value does not match at clock 325");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 326");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 326");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 326");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 326");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 326");
		`Assert(10'b0101000110, OutCounter, "OutCounter: value does not match at clock 326");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 327");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 327");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 327");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 327");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 327");
		`Assert(10'b0101000111, OutCounter, "OutCounter: value does not match at clock 327");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 328");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 328");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 328");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 328");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 328");
		`Assert(10'b0101001000, OutCounter, "OutCounter: value does not match at clock 328");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 329");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 329");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 329");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 329");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 329");
		`Assert(10'b0101001001, OutCounter, "OutCounter: value does not match at clock 329");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 330");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 330");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 330");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 330");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 330");
		`Assert(10'b0101001010, OutCounter, "OutCounter: value does not match at clock 330");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 331");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 331");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 331");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 331");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 331");
		`Assert(10'b0101001011, OutCounter, "OutCounter: value does not match at clock 331");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 332");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 332");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 332");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 332");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 332");
		`Assert(10'b0101001100, OutCounter, "OutCounter: value does not match at clock 332");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 333");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 333");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 333");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 333");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 333");
		`Assert(10'b0101001101, OutCounter, "OutCounter: value does not match at clock 333");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 334");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 334");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 334");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 334");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 334");
		`Assert(10'b0101001110, OutCounter, "OutCounter: value does not match at clock 334");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 335");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 335");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 335");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 335");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 335");
		`Assert(10'b0101001111, OutCounter, "OutCounter: value does not match at clock 335");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 336");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 336");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 336");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 336");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 336");
		`Assert(10'b0101010000, OutCounter, "OutCounter: value does not match at clock 336");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 337");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 337");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 337");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 337");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 337");
		`Assert(10'b0101010001, OutCounter, "OutCounter: value does not match at clock 337");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 338");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 338");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 338");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 338");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 338");
		`Assert(10'b0101010010, OutCounter, "OutCounter: value does not match at clock 338");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 339");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 339");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 339");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 339");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 339");
		`Assert(10'b0101010011, OutCounter, "OutCounter: value does not match at clock 339");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 340");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 340");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 340");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 340");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 340");
		`Assert(10'b0101010100, OutCounter, "OutCounter: value does not match at clock 340");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 341");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 341");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 341");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 341");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 341");
		`Assert(10'b0101010101, OutCounter, "OutCounter: value does not match at clock 341");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 342");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 342");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 342");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 342");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 342");
		`Assert(10'b0101010110, OutCounter, "OutCounter: value does not match at clock 342");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 343");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 343");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 343");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 343");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 343");
		`Assert(10'b0101010111, OutCounter, "OutCounter: value does not match at clock 343");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 344");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 344");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 344");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 344");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 344");
		`Assert(10'b0101011000, OutCounter, "OutCounter: value does not match at clock 344");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 345");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 345");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 345");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 345");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 345");
		`Assert(10'b0101011001, OutCounter, "OutCounter: value does not match at clock 345");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 346");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 346");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 346");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 346");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 346");
		`Assert(10'b0101011010, OutCounter, "OutCounter: value does not match at clock 346");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 347");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 347");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 347");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 347");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 347");
		`Assert(10'b0101011011, OutCounter, "OutCounter: value does not match at clock 347");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 348");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 348");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 348");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 348");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 348");
		`Assert(10'b0101011100, OutCounter, "OutCounter: value does not match at clock 348");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 349");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 349");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 349");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 349");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 349");
		`Assert(10'b0101011101, OutCounter, "OutCounter: value does not match at clock 349");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 350");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 350");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 350");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 350");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 350");
		`Assert(10'b0101011110, OutCounter, "OutCounter: value does not match at clock 350");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 351");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 351");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 351");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 351");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 351");
		`Assert(10'b0101011111, OutCounter, "OutCounter: value does not match at clock 351");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 352");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 352");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 352");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 352");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 352");
		`Assert(10'b0101100000, OutCounter, "OutCounter: value does not match at clock 352");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 353");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 353");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 353");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 353");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 353");
		`Assert(10'b0101100001, OutCounter, "OutCounter: value does not match at clock 353");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 354");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 354");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 354");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 354");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 354");
		`Assert(10'b0101100010, OutCounter, "OutCounter: value does not match at clock 354");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 355");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 355");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 355");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 355");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 355");
		`Assert(10'b0101100011, OutCounter, "OutCounter: value does not match at clock 355");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 356");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 356");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 356");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 356");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 356");
		`Assert(10'b0101100100, OutCounter, "OutCounter: value does not match at clock 356");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 357");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 357");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 357");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 357");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 357");
		`Assert(10'b0101100101, OutCounter, "OutCounter: value does not match at clock 357");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 358");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 358");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 358");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 358");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 358");
		`Assert(10'b0101100110, OutCounter, "OutCounter: value does not match at clock 358");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 359");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 359");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 359");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 359");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 359");
		`Assert(10'b0101100111, OutCounter, "OutCounter: value does not match at clock 359");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 360");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 360");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 360");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 360");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 360");
		`Assert(10'b0101101000, OutCounter, "OutCounter: value does not match at clock 360");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 361");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 361");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 361");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 361");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 361");
		`Assert(10'b0101101001, OutCounter, "OutCounter: value does not match at clock 361");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 362");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 362");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 362");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 362");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 362");
		`Assert(10'b0101101010, OutCounter, "OutCounter: value does not match at clock 362");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 363");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 363");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 363");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 363");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 363");
		`Assert(10'b0101101011, OutCounter, "OutCounter: value does not match at clock 363");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 364");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 364");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 364");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 364");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 364");
		`Assert(10'b0101101100, OutCounter, "OutCounter: value does not match at clock 364");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 365");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 365");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 365");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 365");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 365");
		`Assert(10'b0101101101, OutCounter, "OutCounter: value does not match at clock 365");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 366");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 366");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 366");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 366");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 366");
		`Assert(10'b0101101110, OutCounter, "OutCounter: value does not match at clock 366");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 367");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 367");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 367");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 367");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 367");
		`Assert(10'b0101101111, OutCounter, "OutCounter: value does not match at clock 367");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 368");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 368");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 368");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 368");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 368");
		`Assert(10'b0101110000, OutCounter, "OutCounter: value does not match at clock 368");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 369");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 369");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 369");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 369");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 369");
		`Assert(10'b0101110001, OutCounter, "OutCounter: value does not match at clock 369");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 370");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 370");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 370");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 370");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 370");
		`Assert(10'b0101110010, OutCounter, "OutCounter: value does not match at clock 370");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 371");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 371");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 371");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 371");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 371");
		`Assert(10'b0101110011, OutCounter, "OutCounter: value does not match at clock 371");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 372");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 372");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 372");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 372");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 372");
		`Assert(10'b0101110100, OutCounter, "OutCounter: value does not match at clock 372");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 373");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 373");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 373");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 373");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 373");
		`Assert(10'b0101110101, OutCounter, "OutCounter: value does not match at clock 373");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 374");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 374");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 374");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 374");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 374");
		`Assert(10'b0101110110, OutCounter, "OutCounter: value does not match at clock 374");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 375");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 375");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 375");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 375");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 375");
		`Assert(10'b0101110111, OutCounter, "OutCounter: value does not match at clock 375");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 376");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 376");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 376");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 376");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 376");
		`Assert(10'b0101111000, OutCounter, "OutCounter: value does not match at clock 376");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 377");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 377");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 377");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 377");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 377");
		`Assert(10'b0101111001, OutCounter, "OutCounter: value does not match at clock 377");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 378");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 378");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 378");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 378");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 378");
		`Assert(10'b0101111010, OutCounter, "OutCounter: value does not match at clock 378");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 379");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 379");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 379");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 379");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 379");
		`Assert(10'b0101111011, OutCounter, "OutCounter: value does not match at clock 379");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 380");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 380");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 380");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 380");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 380");
		`Assert(10'b0101111100, OutCounter, "OutCounter: value does not match at clock 380");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 381");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 381");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 381");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 381");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 381");
		`Assert(10'b0101111101, OutCounter, "OutCounter: value does not match at clock 381");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 382");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 382");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 382");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 382");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 382");
		`Assert(10'b0101111110, OutCounter, "OutCounter: value does not match at clock 382");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 383");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 383");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 383");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 383");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 383");
		`Assert(10'b0101111111, OutCounter, "OutCounter: value does not match at clock 383");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 384");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 384");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 384");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 384");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 384");
		`Assert(10'b0110000000, OutCounter, "OutCounter: value does not match at clock 384");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 385");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 385");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 385");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 385");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 385");
		`Assert(10'b0110000001, OutCounter, "OutCounter: value does not match at clock 385");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 386");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 386");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 386");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 386");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 386");
		`Assert(10'b0110000010, OutCounter, "OutCounter: value does not match at clock 386");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 387");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 387");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 387");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 387");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 387");
		`Assert(10'b0110000011, OutCounter, "OutCounter: value does not match at clock 387");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 388");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 388");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 388");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 388");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 388");
		`Assert(10'b0110000100, OutCounter, "OutCounter: value does not match at clock 388");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 389");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 389");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 389");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 389");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 389");
		`Assert(10'b0110000101, OutCounter, "OutCounter: value does not match at clock 389");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 390");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 390");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 390");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 390");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 390");
		`Assert(10'b0110000110, OutCounter, "OutCounter: value does not match at clock 390");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 391");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 391");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 391");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 391");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 391");
		`Assert(10'b0110000111, OutCounter, "OutCounter: value does not match at clock 391");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 392");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 392");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 392");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 392");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 392");
		`Assert(10'b0110001000, OutCounter, "OutCounter: value does not match at clock 392");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 393");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 393");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 393");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 393");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 393");
		`Assert(10'b0110001001, OutCounter, "OutCounter: value does not match at clock 393");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 394");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 394");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 394");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 394");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 394");
		`Assert(10'b0110001010, OutCounter, "OutCounter: value does not match at clock 394");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 395");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 395");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 395");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 395");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 395");
		`Assert(10'b0110001011, OutCounter, "OutCounter: value does not match at clock 395");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 396");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 396");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 396");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 396");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 396");
		`Assert(10'b0110001100, OutCounter, "OutCounter: value does not match at clock 396");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 397");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 397");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 397");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 397");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 397");
		`Assert(10'b0110001101, OutCounter, "OutCounter: value does not match at clock 397");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 398");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 398");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 398");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 398");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 398");
		`Assert(10'b0110001110, OutCounter, "OutCounter: value does not match at clock 398");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 399");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 399");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 399");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 399");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 399");
		`Assert(10'b0110001111, OutCounter, "OutCounter: value does not match at clock 399");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 400");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 400");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 400");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 400");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 400");
		`Assert(10'b0110010000, OutCounter, "OutCounter: value does not match at clock 400");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 401");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 401");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 401");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 401");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 401");
		`Assert(10'b0110010001, OutCounter, "OutCounter: value does not match at clock 401");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 402");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 402");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 402");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 402");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 402");
		`Assert(10'b0110010010, OutCounter, "OutCounter: value does not match at clock 402");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 403");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 403");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 403");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 403");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 403");
		`Assert(10'b0110010011, OutCounter, "OutCounter: value does not match at clock 403");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 404");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 404");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 404");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 404");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 404");
		`Assert(10'b0110010100, OutCounter, "OutCounter: value does not match at clock 404");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 405");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 405");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 405");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 405");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 405");
		`Assert(10'b0110010101, OutCounter, "OutCounter: value does not match at clock 405");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 406");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 406");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 406");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 406");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 406");
		`Assert(10'b0110010110, OutCounter, "OutCounter: value does not match at clock 406");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 407");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 407");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 407");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 407");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 407");
		`Assert(10'b0110010111, OutCounter, "OutCounter: value does not match at clock 407");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 408");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 408");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 408");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 408");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 408");
		`Assert(10'b0110011000, OutCounter, "OutCounter: value does not match at clock 408");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 409");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 409");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 409");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 409");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 409");
		`Assert(10'b0110011001, OutCounter, "OutCounter: value does not match at clock 409");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 410");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 410");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 410");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 410");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 410");
		`Assert(10'b0110011010, OutCounter, "OutCounter: value does not match at clock 410");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 411");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 411");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 411");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 411");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 411");
		`Assert(10'b0110011011, OutCounter, "OutCounter: value does not match at clock 411");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 412");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 412");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 412");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 412");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 412");
		`Assert(10'b0110011100, OutCounter, "OutCounter: value does not match at clock 412");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 413");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 413");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 413");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 413");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 413");
		`Assert(10'b0110011101, OutCounter, "OutCounter: value does not match at clock 413");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 414");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 414");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 414");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 414");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 414");
		`Assert(10'b0110011110, OutCounter, "OutCounter: value does not match at clock 414");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 415");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 415");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 415");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 415");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 415");
		`Assert(10'b0110011111, OutCounter, "OutCounter: value does not match at clock 415");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 416");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 416");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 416");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 416");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 416");
		`Assert(10'b0110100000, OutCounter, "OutCounter: value does not match at clock 416");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 417");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 417");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 417");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 417");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 417");
		`Assert(10'b0110100001, OutCounter, "OutCounter: value does not match at clock 417");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 418");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 418");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 418");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 418");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 418");
		`Assert(10'b0110100010, OutCounter, "OutCounter: value does not match at clock 418");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 419");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 419");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 419");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 419");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 419");
		`Assert(10'b0110100011, OutCounter, "OutCounter: value does not match at clock 419");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 420");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 420");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 420");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 420");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 420");
		`Assert(10'b0110100100, OutCounter, "OutCounter: value does not match at clock 420");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 421");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 421");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 421");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 421");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 421");
		`Assert(10'b0110100101, OutCounter, "OutCounter: value does not match at clock 421");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 422");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 422");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 422");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 422");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 422");
		`Assert(10'b0110100110, OutCounter, "OutCounter: value does not match at clock 422");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 423");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 423");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 423");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 423");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 423");
		`Assert(10'b0110100111, OutCounter, "OutCounter: value does not match at clock 423");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 424");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 424");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 424");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 424");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 424");
		`Assert(10'b0110101000, OutCounter, "OutCounter: value does not match at clock 424");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 425");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 425");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 425");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 425");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 425");
		`Assert(10'b0110101001, OutCounter, "OutCounter: value does not match at clock 425");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 426");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 426");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 426");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 426");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 426");
		`Assert(10'b0110101010, OutCounter, "OutCounter: value does not match at clock 426");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 427");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 427");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 427");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 427");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 427");
		`Assert(10'b0110101011, OutCounter, "OutCounter: value does not match at clock 427");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 428");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 428");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 428");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 428");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 428");
		`Assert(10'b0110101100, OutCounter, "OutCounter: value does not match at clock 428");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 429");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 429");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 429");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 429");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 429");
		`Assert(10'b0110101101, OutCounter, "OutCounter: value does not match at clock 429");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 430");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 430");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 430");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 430");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 430");
		`Assert(10'b0110101110, OutCounter, "OutCounter: value does not match at clock 430");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 431");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 431");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 431");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 431");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 431");
		`Assert(10'b0110101111, OutCounter, "OutCounter: value does not match at clock 431");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 432");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 432");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 432");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 432");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 432");
		`Assert(10'b0110110000, OutCounter, "OutCounter: value does not match at clock 432");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 433");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 433");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 433");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 433");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 433");
		`Assert(10'b0110110001, OutCounter, "OutCounter: value does not match at clock 433");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 434");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 434");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 434");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 434");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 434");
		`Assert(10'b0110110010, OutCounter, "OutCounter: value does not match at clock 434");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 435");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 435");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 435");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 435");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 435");
		`Assert(10'b0110110011, OutCounter, "OutCounter: value does not match at clock 435");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 436");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 436");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 436");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 436");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 436");
		`Assert(10'b0110110100, OutCounter, "OutCounter: value does not match at clock 436");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 437");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 437");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 437");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 437");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 437");
		`Assert(10'b0110110101, OutCounter, "OutCounter: value does not match at clock 437");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 438");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 438");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 438");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 438");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 438");
		`Assert(10'b0110110110, OutCounter, "OutCounter: value does not match at clock 438");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 439");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 439");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 439");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 439");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 439");
		`Assert(10'b0110110111, OutCounter, "OutCounter: value does not match at clock 439");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 440");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 440");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 440");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 440");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 440");
		`Assert(10'b0110111000, OutCounter, "OutCounter: value does not match at clock 440");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 441");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 441");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 441");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 441");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 441");
		`Assert(10'b0110111001, OutCounter, "OutCounter: value does not match at clock 441");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 442");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 442");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 442");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 442");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 442");
		`Assert(10'b0110111010, OutCounter, "OutCounter: value does not match at clock 442");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 443");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 443");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 443");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 443");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 443");
		`Assert(10'b0110111011, OutCounter, "OutCounter: value does not match at clock 443");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 444");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 444");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 444");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 444");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 444");
		`Assert(10'b0110111100, OutCounter, "OutCounter: value does not match at clock 444");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 445");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 445");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 445");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 445");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 445");
		`Assert(10'b0110111101, OutCounter, "OutCounter: value does not match at clock 445");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 446");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 446");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 446");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 446");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 446");
		`Assert(10'b0110111110, OutCounter, "OutCounter: value does not match at clock 446");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 447");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 447");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 447");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 447");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 447");
		`Assert(10'b0110111111, OutCounter, "OutCounter: value does not match at clock 447");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 448");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 448");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 448");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 448");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 448");
		`Assert(10'b0111000000, OutCounter, "OutCounter: value does not match at clock 448");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 449");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 449");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 449");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 449");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 449");
		`Assert(10'b0111000001, OutCounter, "OutCounter: value does not match at clock 449");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 450");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 450");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 450");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 450");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 450");
		`Assert(10'b0111000010, OutCounter, "OutCounter: value does not match at clock 450");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 451");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 451");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 451");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 451");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 451");
		`Assert(10'b0111000011, OutCounter, "OutCounter: value does not match at clock 451");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 452");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 452");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 452");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 452");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 452");
		`Assert(10'b0111000100, OutCounter, "OutCounter: value does not match at clock 452");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 453");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 453");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 453");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 453");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 453");
		`Assert(10'b0111000101, OutCounter, "OutCounter: value does not match at clock 453");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 454");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 454");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 454");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 454");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 454");
		`Assert(10'b0111000110, OutCounter, "OutCounter: value does not match at clock 454");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 455");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 455");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 455");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 455");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 455");
		`Assert(10'b0111000111, OutCounter, "OutCounter: value does not match at clock 455");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 456");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 456");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 456");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 456");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 456");
		`Assert(10'b0111001000, OutCounter, "OutCounter: value does not match at clock 456");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 457");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 457");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 457");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 457");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 457");
		`Assert(10'b0111001001, OutCounter, "OutCounter: value does not match at clock 457");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 458");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 458");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 458");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 458");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 458");
		`Assert(10'b0111001010, OutCounter, "OutCounter: value does not match at clock 458");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 459");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 459");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 459");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 459");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 459");
		`Assert(10'b0111001011, OutCounter, "OutCounter: value does not match at clock 459");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 460");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 460");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 460");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 460");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 460");
		`Assert(10'b0111001100, OutCounter, "OutCounter: value does not match at clock 460");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 461");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 461");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 461");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 461");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 461");
		`Assert(10'b0111001101, OutCounter, "OutCounter: value does not match at clock 461");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 462");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 462");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 462");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 462");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 462");
		`Assert(10'b0111001110, OutCounter, "OutCounter: value does not match at clock 462");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 463");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 463");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 463");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 463");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 463");
		`Assert(10'b0111001111, OutCounter, "OutCounter: value does not match at clock 463");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 464");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 464");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 464");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 464");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 464");
		`Assert(10'b0111010000, OutCounter, "OutCounter: value does not match at clock 464");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 465");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 465");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 465");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 465");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 465");
		`Assert(10'b0111010001, OutCounter, "OutCounter: value does not match at clock 465");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 466");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 466");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 466");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 466");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 466");
		`Assert(10'b0111010010, OutCounter, "OutCounter: value does not match at clock 466");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 467");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 467");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 467");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 467");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 467");
		`Assert(10'b0111010011, OutCounter, "OutCounter: value does not match at clock 467");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 468");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 468");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 468");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 468");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 468");
		`Assert(10'b0111010100, OutCounter, "OutCounter: value does not match at clock 468");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 469");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 469");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 469");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 469");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 469");
		`Assert(10'b0111010101, OutCounter, "OutCounter: value does not match at clock 469");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 470");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 470");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 470");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 470");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 470");
		`Assert(10'b0111010110, OutCounter, "OutCounter: value does not match at clock 470");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 471");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 471");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 471");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 471");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 471");
		`Assert(10'b0111010111, OutCounter, "OutCounter: value does not match at clock 471");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 472");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 472");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 472");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 472");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 472");
		`Assert(10'b0111011000, OutCounter, "OutCounter: value does not match at clock 472");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 473");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 473");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 473");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 473");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 473");
		`Assert(10'b0111011001, OutCounter, "OutCounter: value does not match at clock 473");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 474");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 474");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 474");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 474");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 474");
		`Assert(10'b0111011010, OutCounter, "OutCounter: value does not match at clock 474");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 475");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 475");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 475");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 475");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 475");
		`Assert(10'b0111011011, OutCounter, "OutCounter: value does not match at clock 475");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 476");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 476");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 476");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 476");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 476");
		`Assert(10'b0111011100, OutCounter, "OutCounter: value does not match at clock 476");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 477");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 477");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 477");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 477");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 477");
		`Assert(10'b0111011101, OutCounter, "OutCounter: value does not match at clock 477");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 478");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 478");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 478");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 478");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 478");
		`Assert(10'b0111011110, OutCounter, "OutCounter: value does not match at clock 478");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 479");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 479");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 479");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 479");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 479");
		`Assert(10'b0111011111, OutCounter, "OutCounter: value does not match at clock 479");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 480");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 480");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 480");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 480");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 480");
		`Assert(10'b0111100000, OutCounter, "OutCounter: value does not match at clock 480");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 481");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 481");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 481");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 481");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 481");
		`Assert(10'b0111100001, OutCounter, "OutCounter: value does not match at clock 481");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 482");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 482");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 482");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 482");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 482");
		`Assert(10'b0111100010, OutCounter, "OutCounter: value does not match at clock 482");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 483");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 483");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 483");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 483");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 483");
		`Assert(10'b0111100011, OutCounter, "OutCounter: value does not match at clock 483");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 484");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 484");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 484");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 484");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 484");
		`Assert(10'b0111100100, OutCounter, "OutCounter: value does not match at clock 484");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 485");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 485");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 485");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 485");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 485");
		`Assert(10'b0111100101, OutCounter, "OutCounter: value does not match at clock 485");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 486");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 486");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 486");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 486");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 486");
		`Assert(10'b0111100110, OutCounter, "OutCounter: value does not match at clock 486");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 487");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 487");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 487");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 487");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 487");
		`Assert(10'b0111100111, OutCounter, "OutCounter: value does not match at clock 487");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 488");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 488");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 488");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 488");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 488");
		`Assert(10'b0111101000, OutCounter, "OutCounter: value does not match at clock 488");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 489");
		`Assert(1'b1, OutFP, "OutFP: value does not match at clock 489");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 489");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 489");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 489");
		`Assert(10'b0111101001, OutCounter, "OutCounter: value does not match at clock 489");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 490");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 490");
		`Assert(1'b1, OutSP, "OutSP: value does not match at clock 490");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 490");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 490");
		`Assert(10'b0111101010, OutCounter, "OutCounter: value does not match at clock 490");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 491");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 491");
		`Assert(1'b1, OutSP, "OutSP: value does not match at clock 491");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 491");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 491");
		`Assert(10'b0111101011, OutCounter, "OutCounter: value does not match at clock 491");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 492");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 492");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 492");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 492");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 492");
		`Assert(10'b0111101100, OutCounter, "OutCounter: value does not match at clock 492");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 493");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 493");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 493");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 493");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 493");
		`Assert(10'b0111101101, OutCounter, "OutCounter: value does not match at clock 493");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 494");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 494");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 494");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 494");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 494");
		`Assert(10'b0111101110, OutCounter, "OutCounter: value does not match at clock 494");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 495");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 495");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 495");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 495");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 495");
		`Assert(10'b0111101111, OutCounter, "OutCounter: value does not match at clock 495");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 496");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 496");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 496");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 496");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 496");
		`Assert(10'b0111110000, OutCounter, "OutCounter: value does not match at clock 496");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 497");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 497");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 497");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 497");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 497");
		`Assert(10'b0111110001, OutCounter, "OutCounter: value does not match at clock 497");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 498");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 498");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 498");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 498");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 498");
		`Assert(10'b0111110010, OutCounter, "OutCounter: value does not match at clock 498");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 499");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 499");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 499");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 499");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 499");
		`Assert(10'b0111110011, OutCounter, "OutCounter: value does not match at clock 499");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 500");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 500");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 500");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 500");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 500");
		`Assert(10'b0111110100, OutCounter, "OutCounter: value does not match at clock 500");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 501");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 501");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 501");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 501");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 501");
		`Assert(10'b0111110101, OutCounter, "OutCounter: value does not match at clock 501");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 502");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 502");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 502");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 502");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 502");
		`Assert(10'b0111110110, OutCounter, "OutCounter: value does not match at clock 502");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 503");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 503");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 503");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 503");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 503");
		`Assert(10'b0111110111, OutCounter, "OutCounter: value does not match at clock 503");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 504");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 504");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 504");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 504");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 504");
		`Assert(10'b0111111000, OutCounter, "OutCounter: value does not match at clock 504");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 505");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 505");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 505");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 505");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 505");
		`Assert(10'b0111111001, OutCounter, "OutCounter: value does not match at clock 505");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 506");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 506");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 506");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 506");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 506");
		`Assert(10'b0111111010, OutCounter, "OutCounter: value does not match at clock 506");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 507");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 507");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 507");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 507");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 507");
		`Assert(10'b0111111011, OutCounter, "OutCounter: value does not match at clock 507");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 508");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 508");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 508");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 508");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 508");
		`Assert(10'b0111111100, OutCounter, "OutCounter: value does not match at clock 508");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 509");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 509");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 509");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 509");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 509");
		`Assert(10'b0111111101, OutCounter, "OutCounter: value does not match at clock 509");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 510");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 510");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 510");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 510");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 510");
		`Assert(10'b0111111110, OutCounter, "OutCounter: value does not match at clock 510");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 511");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 511");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 511");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 511");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 511");
		`Assert(10'b0111111111, OutCounter, "OutCounter: value does not match at clock 511");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 512");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 512");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 512");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 512");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 512");
		`Assert(10'b1000000000, OutCounter, "OutCounter: value does not match at clock 512");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 513");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 513");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 513");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 513");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 513");
		`Assert(10'b1000000001, OutCounter, "OutCounter: value does not match at clock 513");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 514");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 514");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 514");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 514");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 514");
		`Assert(10'b1000000010, OutCounter, "OutCounter: value does not match at clock 514");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 515");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 515");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 515");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 515");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 515");
		`Assert(10'b1000000011, OutCounter, "OutCounter: value does not match at clock 515");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 516");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 516");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 516");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 516");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 516");
		`Assert(10'b1000000100, OutCounter, "OutCounter: value does not match at clock 516");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 517");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 517");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 517");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 517");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 517");
		`Assert(10'b1000000101, OutCounter, "OutCounter: value does not match at clock 517");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 518");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 518");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 518");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 518");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 518");
		`Assert(10'b1000000110, OutCounter, "OutCounter: value does not match at clock 518");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 519");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 519");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 519");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 519");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 519");
		`Assert(10'b1000000111, OutCounter, "OutCounter: value does not match at clock 519");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 520");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 520");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 520");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 520");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 520");
		`Assert(10'b1000001000, OutCounter, "OutCounter: value does not match at clock 520");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 521");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 521");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 521");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 521");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 521");
		`Assert(10'b1000001001, OutCounter, "OutCounter: value does not match at clock 521");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 522");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 522");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 522");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 522");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 522");
		`Assert(10'b1000001010, OutCounter, "OutCounter: value does not match at clock 522");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 523");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 523");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 523");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 523");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 523");
		`Assert(10'b1000001011, OutCounter, "OutCounter: value does not match at clock 523");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b0, OutVisible, "OutVisible: value does not match at clock 524");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 524");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 524");
		`Assert(1'b1, OutBP, "OutBP: value does not match at clock 524");
		`Assert(1'b1, OutMax, "OutMax: value does not match at clock 524");
		`Assert(10'b1000001100, OutCounter, "OutCounter: value does not match at clock 524");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 525");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 525");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 525");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 525");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 525");
		`Assert(10'b0000000000, OutCounter, "OutCounter: value does not match at clock 525");

		Enabled = 1'b1;
		@(negedge clk);
		`Assert(1'b1, OutVisible, "OutVisible: value does not match at clock 526");
		`Assert(1'b0, OutFP, "OutFP: value does not match at clock 526");
		`Assert(1'b0, OutSP, "OutSP: value does not match at clock 526");
		`Assert(1'b0, OutBP, "OutBP: value does not match at clock 526");
		`Assert(1'b0, OutMax, "OutMax: value does not match at clock 526");
		`Assert(10'b0000000001, OutCounter, "OutCounter: value does not match at clock 526");
	end

	// DUT instantiation
	VGASyncModule_TopLevel dut (
		.Clock (clk),
		.Reset (reset),
		.Enabled (Enabled),
		.OutVisible (OutVisible),
		.OutFP (OutFP),
		.OutSP (OutSP),
		.OutBP (OutBP),
		.OutMax (OutMax),
		.OutCounter (OutCounter)
	);
endmodule
